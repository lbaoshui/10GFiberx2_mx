library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity vsync_cross is
generic
(
    DLY_CY : integer := 3
);
port 
(
    vsync_async     : in std_logic; 
    nRST            : in std_logic;
    clk             : in std_logic; 
    vsync_synced    : out std_logic 
);
end vsync_cross;

architecture behaviour of vsync_cross is
 
signal vsync_buf_sys        : std_logic_vector(DLY_CY-1 downto 0) := (others=>'0');
signal vsync_final          : std_logic :='0';

begin 

process(nRST,clk)
begin
    if nRST = '0' then
        vsync_buf_sys <= (OTHERS=>'0');
        vsync_final   <= '0';
    elsif rising_edge(clk) then
        vsync_buf_sys <= vsync_buf_sys(DLY_CY-2 downto 0) & vsync_async;
        vsync_final   <= vsync_buf_sys(DLY_CY-1);
    end if;
end process;

vsync_synced <= vsync_final;

end;