// issp.v

// Generated using ACDS version 21.3 170

`timescale 1 ps / 1 ps
module issp (
		output wire [1:0] source, // sources.source
		input  wire [0:0] probe   //  probes.probe
	);

	altsource_probe #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (1),
		.source_width            (2),
		.source_initial_value    ("0"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.source     (source), //  output,  width = 2, sources.source
		.probe      (probe),  //   input,  width = 1,  probes.probe
		.source_ena (1'b1)    // (terminated),                     
	);

endmodule
