module probe_flow (
		output wire [31:0] source, // sources.source
		input  wire [0:0]  probe   //  probes.probe
	);
endmodule

