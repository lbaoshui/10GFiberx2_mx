module Probe (
		output wire [3:0] source,     //    sources.source
		input  wire       source_clk, // source_clk.clk
		input  wire [0:0] probe       //     probes.probe
	);
endmodule

