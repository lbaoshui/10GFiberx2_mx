library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.PCK_bk_serdes.all;

entity BK2fiber_pack is 

end BK2fiber_pack;

architecture beha of BK2fiber_pack is 

begin 



end beha;