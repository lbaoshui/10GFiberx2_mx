module issp (
		output wire [1:0] source, // sources.source
		input  wire [0:0] probe   //  probes.probe
	);
endmodule

