module LPM_9x10 (
		input  wire [9:0]  dataa,  //  dataa.dataa
		output wire [18:0] result, // result.result
		input  wire [8:0]  datab,  //  datab.datab
		input  wire        clock   //  clock.clk
	);
endmodule

