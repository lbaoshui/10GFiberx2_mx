-- generic_spi_flash.vhd

-- Generated using ACDS version 18.1 222

library IEEE;
library intel_generic_serial_flash_interface_top_181;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity generic_spi_flash is
	port (
		avl_csr_address       : in  std_logic_vector(5 downto 0)  := (others => '0'); -- avl_csr.address
		avl_csr_read          : in  std_logic                     := '0';             --        .read
		avl_csr_readdata      : out std_logic_vector(31 downto 0);                    --        .readdata
		avl_csr_write         : in  std_logic                     := '0';             --        .write
		avl_csr_writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --        .writedata
		avl_csr_waitrequest   : out std_logic;                                        --        .waitrequest
		avl_csr_readdatavalid : out std_logic;                                        --        .readdatavalid
		avl_mem_write         : in  std_logic                     := '0';             -- avl_mem.write
		avl_mem_burstcount    : in  std_logic_vector(6 downto 0)  := (others => '0'); --        .burstcount
		avl_mem_waitrequest   : out std_logic;                                        --        .waitrequest
		avl_mem_read          : in  std_logic                     := '0';             --        .read
		avl_mem_address       : in  std_logic_vector(22 downto 0) := (others => '0'); --        .address
		avl_mem_writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --        .writedata
		avl_mem_readdata      : out std_logic_vector(31 downto 0);                    --        .readdata
		avl_mem_readdatavalid : out std_logic;                                        --        .readdatavalid
		avl_mem_byteenable    : in  std_logic_vector(3 downto 0)  := (others => '0'); --        .byteenable
		clk_clk               : in  std_logic                     := '0';             --     clk.clk
		reset_reset           : in  std_logic                     := '0'              --   reset.reset
	);
end entity generic_spi_flash;

architecture rtl of generic_spi_flash is
	component generic_spi_flash_intel_generic_serial_flash_interface_top_181_zqmrk7a_cmp is
		generic (
			DEVICE_FAMILY : string  := "";
			CHIP_SELS     : integer := 1
		);
		port (
			avl_csr_address       : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			avl_csr_read          : in  std_logic                     := 'X';             -- read
			avl_csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avl_csr_write         : in  std_logic                     := 'X';             -- write
			avl_csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_csr_waitrequest   : out std_logic;                                        -- waitrequest
			avl_csr_readdatavalid : out std_logic;                                        -- readdatavalid
			avl_mem_write         : in  std_logic                     := 'X';             -- write
			avl_mem_burstcount    : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			avl_mem_waitrequest   : out std_logic;                                        -- waitrequest
			avl_mem_read          : in  std_logic                     := 'X';             -- read
			avl_mem_address       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			avl_mem_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_mem_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avl_mem_readdatavalid : out std_logic;                                        -- readdatavalid
			avl_mem_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk_clk               : in  std_logic                     := 'X';             -- clk
			reset_reset           : in  std_logic                     := 'X'              -- reset
		);
	end component generic_spi_flash_intel_generic_serial_flash_interface_top_181_zqmrk7a_cmp;

	for intel_generic_serial_flash_interface_top_0 : generic_spi_flash_intel_generic_serial_flash_interface_top_181_zqmrk7a_cmp
		use entity intel_generic_serial_flash_interface_top_181.generic_spi_flash_intel_generic_serial_flash_interface_top_181_zqmrk7a;
begin

	intel_generic_serial_flash_interface_top_0 : component generic_spi_flash_intel_generic_serial_flash_interface_top_181_zqmrk7a_cmp
		generic map (
			DEVICE_FAMILY => "Arria 10",
			CHIP_SELS     => 1
		)
		port map (
			avl_csr_address       => avl_csr_address,       -- avl_csr.address
			avl_csr_read          => avl_csr_read,          --        .read
			avl_csr_readdata      => avl_csr_readdata,      --        .readdata
			avl_csr_write         => avl_csr_write,         --        .write
			avl_csr_writedata     => avl_csr_writedata,     --        .writedata
			avl_csr_waitrequest   => avl_csr_waitrequest,   --        .waitrequest
			avl_csr_readdatavalid => avl_csr_readdatavalid, --        .readdatavalid
			avl_mem_write         => avl_mem_write,         -- avl_mem.write
			avl_mem_burstcount    => avl_mem_burstcount,    --        .burstcount
			avl_mem_waitrequest   => avl_mem_waitrequest,   --        .waitrequest
			avl_mem_read          => avl_mem_read,          --        .read
			avl_mem_address       => avl_mem_address,       --        .address
			avl_mem_writedata     => avl_mem_writedata,     --        .writedata
			avl_mem_readdata      => avl_mem_readdata,      --        .readdata
			avl_mem_readdatavalid => avl_mem_readdatavalid, --        .readdatavalid
			avl_mem_byteenable    => avl_mem_byteenable,    --        .byteenable
			clk_clk               => clk_clk,               --     clk.clk
			reset_reset           => reset_reset            --   reset.reset
		);

end architecture rtl; -- of generic_spi_flash
