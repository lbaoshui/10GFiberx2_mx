library IEEE;
use IEEE.std_logic_1164.all;
--PCK_version for 027 FPGA .
package PCK_version_FPGA_def is

constant     PCK_CONS_VER_HIGH           : std_logic_vector  :=X"03";
constant     PCK_CONS_VER_LOW            : std_logic_vector  :=X"04";
constant     PCK_PCB_M_VER               : std_logic_vector  :=x"01"; --NOT USED 
constant     PCK_PCB_S_VER               : std_logic_vector  :=X"00"; --NOT USED 

--0: 027
--1: 032 
constant     FPGA032_EN             : integer := 0;   --20221122 wangac 
 
end PCK_version_FPGA_def;

library IEEE;
use IEEE.std_logic_1164.all;

package body PCK_version_FPGA_def is


end PCK_version_FPGA_def;