// fifo320.v

// Generated using ACDS version 18.1 222

`timescale 1 ps / 1 ps
module fifo320 (
		input  wire [319:0] data,  //  fifo_input.datain
		input  wire         wrreq, //            .wrreq
		input  wire         rdreq, //            .rdreq
		input  wire         clock, //            .clk
		input  wire         aclr,  //            .aclr
		output wire [319:0] q,     // fifo_output.dataout
		output wire         full,  //            .full
		output wire         empty  //            .empty
	);

	fifo320_fifo_181_hlc74wy fifo_0 (
		.data  (data),  //   input,  width = 320,  fifo_input.datain
		.wrreq (wrreq), //   input,    width = 1,            .wrreq
		.rdreq (rdreq), //   input,    width = 1,            .rdreq
		.clock (clock), //   input,    width = 1,            .clk
		.aclr  (aclr),  //   input,    width = 1,            .aclr
		.q     (q),     //  output,  width = 320, fifo_output.dataout
		.full  (full),  //  output,    width = 1,            .full
		.empty (empty)  //  output,    width = 1,            .empty
	);

endmodule
